package AES;

import AES_Defs :: *;
export AES_Defs :: *;

import AES_Encrypt_Decrypt :: *;
export AES_Encrypt_Decrypt :: *;

import AES_IFCs :: *;
export AES_IFCs :: *;

import AES_KeyExpand :: *;
export AES_KeyExpand :: *;

import AES_Params :: *;
export AES_Params :: *;

endpackage